module uart_rx #(
    parameter int BAUD_DIV = 434,  // BAUD_DIV = 50M / 115200 ≈ 434
    // cứ 434clk thì gửi 1 bit, chia 434clk ra thành 27tick, mỗi tick lấy mẫu data 1 lần
    parameter int TICK_DIV = 27    // số chu kỳ clock mỗi tick (~27)
                                   // tick_div = Ttick/Tclk (Ttick = Tbit/16sampling)
)(
    input  logic clk,              // Xung clock 50 MHz
    input  logic rst_n,            // Reset active-low
    input  logic rx,               // Đầu vào UART RX
    output logic [7:0] data_out,   // Dữ liệu nhận được
    output logic valid             // Báo hiệu dữ liệu hợp lệ
);
    // --- State encoding
    localparam int STATE_IDLE  = 2'd0;
    localparam int STATE_START = 2'd1;
    localparam int STATE_DATA  = 2'd2;
    localparam int STATE_STOP  = 2'd3;
    // --- Internal registers
    logic [1:0] state;
    logic [12:0] clk_counter;
    logic [3:0]  tick_counter;
    logic [3:0]  bit_index;
    logic [7:0]  rx_shift;
    logic        rx_sync1, rx_sync2; //Đồng bộ hóa tín hiệu rx
    // --- Đồng bộ hóa tín hiệu RX
	 //
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            rx_sync1 <= 1'b1;
            rx_sync2 <= 1'b1;
        end else begin
            rx_sync1 <= rx;
            rx_sync2 <= rx_sync1;
        end
    end
//

    // --- FSM nhận UART
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state        <= STATE_IDLE;
            clk_counter  <= 13'd0;
            tick_counter <= 4'd0;
            bit_index    <= 4'd0;
            rx_shift     <= 8'd0;
            data_out     <= 8'd0;
            valid        <= 1'b0;
				
        end else begin
            case (state)
                STATE_IDLE: begin
                    valid        <= 1'b0;
                    clk_counter  <= 13'd0;
                    tick_counter <= 4'd0;
                    bit_index    <= 4'd0;

                    if (rx_sync2 == 1'b0) begin
                        state <= STATE_START;
                    end
                end

                STATE_START: begin
                    if (clk_counter < TICK_DIV - 1) begin
                        clk_counter <= clk_counter + 1'b1;
                    end else begin
                        clk_counter  <= 13'd0;
                        tick_counter <= tick_counter + 1'b1;

                        if (tick_counter == 4'd8) begin
                            if (rx_sync2 == 1'b0)
                                state <= STATE_DATA;
                            else
                                state <= STATE_IDLE;
                        end
                    end
                end

                STATE_DATA: begin
                    if (clk_counter < TICK_DIV - 1) begin
                        clk_counter <= clk_counter + 1'b1;
                    end else begin
                        clk_counter  <= 13'd0;
                        tick_counter <= tick_counter + 1'b1;

                        if (tick_counter == 4'd8) begin
                            rx_shift[bit_index] <= rx_sync2;

                            if (bit_index < 4'd7)
                                bit_index <= bit_index + 1'b1;
                            else begin
                                bit_index <= 4'd0;
                                state <= STATE_STOP;
                            end
                        end
                    end
                end

                STATE_STOP: begin
                    if (clk_counter < TICK_DIV - 1) begin
                        clk_counter <= clk_counter + 1'b1;
                    end else begin
                        clk_counter  <= 13'd0;
                        tick_counter <= tick_counter + 1'b1;

                        if (tick_counter == 4'd8) begin
                            if (rx_sync2 == 1'b1) begin
                                data_out <= rx_shift;
                                valid    <= 1'b1;
                            end
                            state <= STATE_IDLE;
                        end
                    end
                end

                
            endcase
        end
    end

endmodule
